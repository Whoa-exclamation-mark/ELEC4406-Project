ENTITY control_unit_tb IS
	
END control_unit_tb;

ARCHITECTURE control_unit_tb_rtl OF control_unit_tb IS

BEGIN

END control_unit_tb_rtl;